library ieee;
use ieee.std_logic_1164.all;

entity bitComparator_tb is
end entity bitComparator_tb;

architecture testbench of bitComparator_tb is
    signal a_tb 		: 	std_logic_vector(3 downto 0) := "0000";
    signal b_tb 		: 	std_logic_vector(3 downto 0) := "0000";
    signal lg_tb 		: 	std_logic;
    signal eq_tb                :       std_logic;
    signal ls_tb                :       std_logic;
begin
    a_tb <=   "0001" after 3200 ns,
	      "0010" after 6400 ns,
	      "0011" after 9600 ns,
              "0100" after 12800 ns,
              "0101" after 16000 ns,
              "0110" after 19200 ns,
              "0111" after 22400 ns,
              "1000" after 25600 ns,
              "1001" after 28800 ns,
              "1010" after 32000 ns,
              "1011" after 35200 ns,
              "1100" after 38400 ns,
              "1101" after 41600 ns,
              "1110" after 44800 ns,
              "1111" after 48000 ns;
    
    b_tb <=   "0001" after 200 ns,
	      "0010" after 400 ns,
	      "0011" after 600 ns,
	      "0100" after 800 ns,
	      "0101" after 1000 ns,
	      "0110" after 1200 ns,
	      "0111" after 1400 ns,
	      "1000" after 1600 ns,
	      "1001" after 1800 ns,
	      "1010" after 2000 ns,
	      "1011" after 2200 ns,
	      "1100" after 2400 ns,
	      "1101" after 2600 ns,
	      "1110" after 2800 ns,
	      "1111" after 3000 ns,
	      --0001
              "0000" after 3200 ns,
	      "0001" after 3400 ns,
	      "0010" after 3600 ns,
	      "0011" after 3800 ns,
	      "0100" after 4000 ns,
	      "0101" after 4200 ns,
	      "0110" after 4400 ns,
	      "0111" after 4600 ns,
	      "1000" after 4800 ns,
	      "1001" after 5000 ns,
	      "1010" after 5200 ns,
	      "1011" after 5400 ns,
	      "1100" after 5600 ns,
	      "1101" after 5800 ns,
	      "1110" after 6000 ns,
	      "1111" after 6200 ns,
              --0010
              "0000" after 6400 ns,
	      "0001" after 6600 ns,
	      "0010" after 6800 ns,
	      "0011" after 7000 ns,
	      "0100" after 7200 ns,
	      "0101" after 7400 ns,
	      "0110" after 7600 ns,
	      "0111" after 7800 ns,
	      "1000" after 8000 ns,
	      "1001" after 8200 ns,
	      "1010" after 8400 ns,
	      "1011" after 8600 ns,
	      "1100" after 8800 ns,
	      "1101" after 9000 ns,
	      "1110" after 9200 ns,
	      "1111" after 9400 ns,
              --0011
              "0000" after 9600 ns,
	      "0001" after 9800 ns,
	      "0010" after 10000 ns,
	      "0011" after 10200 ns,
	      "0100" after 10400 ns,
	      "0101" after 10600 ns,
	      "0110" after 10800 ns,
	      "0111" after 11000 ns,
	      "1000" after 11200 ns,
	      "1001" after 11400 ns,
	      "1010" after 11600 ns,
	      "1011" after 11800 ns,
	      "1100" after 12000 ns,
	      "1101" after 12200 ns,
	      "1110" after 12400 ns,
	      "1111" after 12600 ns,
              --0100
              "0000" after 12800 ns,
	      "0001" after 13000 ns,
	      "0010" after 13200 ns,
	      "0011" after 13400 ns,
	      "0100" after 13600 ns,
	      "0101" after 13800 ns,
	      "0110" after 14000 ns,
	      "0111" after 14200 ns,
	      "1000" after 14400 ns,
	      "1001" after 14600 ns,
	      "1010" after 14800 ns,
	      "1011" after 15000 ns,
	      "1100" after 15200 ns,
	      "1101" after 15400 ns,
	      "1110" after 15600 ns,
	      "1111" after 15800 ns,
              --0101
              "0000" after 16000 ns,
	      "0001" after 16200 ns,
	      "0010" after 16400 ns,
	      "0011" after 16600 ns,
	      "0100" after 16800 ns,
	      "0101" after 17000 ns,
	      "0110" after 17200 ns,
	      "0111" after 17400 ns,
	      "1000" after 17600 ns,
	      "1001" after 17800 ns,
	      "1010" after 18000 ns,
	      "1011" after 18200 ns,
	      "1100" after 18400 ns,
	      "1101" after 18600 ns,
	      "1110" after 18800 ns,
	      "1111" after 19000 ns,
              --0110
              "0000" after 19200 ns,
	      "0001" after 19400 ns,
	      "0010" after 19600 ns,
	      "0011" after 19800 ns,
	      "0100" after 20000 ns,
	      "0101" after 20200 ns,
	      "0110" after 20400 ns,
	      "0111" after 20600 ns,
	      "1000" after 20800 ns,
	      "1001" after 21000 ns,
	      "1010" after 21200 ns,
	      "1011" after 21400 ns,
	      "1100" after 21600 ns,
	      "1101" after 21800 ns,
	      "1110" after 22000 ns,
	      "1111" after 22200 ns,
              --0111
              "0000" after 22400 ns,
	      "0001" after 22600 ns,
	      "0010" after 22800 ns,
	      "0011" after 23000 ns,
	      "0100" after 23200 ns,
	      "0101" after 23400 ns,
	      "0110" after 23600 ns,
	      "0111" after 23800 ns,
	      "1000" after 24000 ns,
	      "1001" after 24200 ns,
	      "1010" after 24400 ns,
	      "1011" after 24600 ns,
	      "1100" after 24800 ns,
	      "1101" after 25000 ns,
	      "1110" after 25200 ns,
	      "1111" after 25400 ns,
              --1000
              "0000" after 25600 ns,
	      "0001" after 25800 ns,
	      "0010" after 26000 ns,
	      "0011" after 26200 ns,
	      "0100" after 26400 ns,
	      "0101" after 26600 ns,
	      "0110" after 26800 ns,
	      "0111" after 27000 ns,
	      "1000" after 27200 ns,
	      "1001" after 27400 ns,
	      "1010" after 27600 ns,
	      "1011" after 27800 ns,
	      "1100" after 28000 ns,
	      "1101" after 28200 ns,
	      "1110" after 28400 ns,
	      "1111" after 28600 ns,
              --1001
              "0000" after 28800 ns,
	      "0001" after 29000 ns,
	      "0010" after 29200 ns,
	      "0011" after 29400 ns,
	      "0100" after 29600 ns,
	      "0101" after 29800 ns,
	      "0110" after 30000 ns,
	      "0111" after 30200 ns,
	      "1000" after 30400 ns,
	      "1001" after 30600 ns,
	      "1010" after 30800 ns,
	      "1011" after 31000 ns,
	      "1100" after 31200 ns,
	      "1101" after 31400 ns,
	      "1110" after 31600 ns,
	      "1111" after 31800 ns,
              --1010
              "0000" after 32000 ns,
	      "0001" after 32200 ns,
	      "0010" after 32400 ns,
	      "0011" after 32600 ns,
	      "0100" after 32800 ns,
	      "0101" after 33000 ns,
	      "0110" after 33200 ns,
	      "0111" after 33400 ns,
	      "1000" after 33600 ns,
	      "1001" after 33800 ns,
	      "1010" after 34000 ns,
	      "1011" after 34200 ns,
	      "1100" after 34400 ns,
	      "1101" after 34600 ns,
	      "1110" after 34800 ns,
	      "1111" after 35000 ns,
              --1011
              "0000" after 35200 ns,
	      "0001" after 35400 ns,
	      "0010" after 35600 ns,
	      "0011" after 35800 ns,
	      "0100" after 36000 ns,
	      "0101" after 36200 ns,
	      "0110" after 36400 ns,
	      "0111" after 36600 ns,
	      "1000" after 36800 ns,
	      "1001" after 37000 ns,
	      "1010" after 37200 ns,
	      "1011" after 37400 ns,
	      "1100" after 37600 ns,
	      "1101" after 37800 ns,
	      "1110" after 38000 ns,
	      "1111" after 38200 ns,
              --1100
              "0000" after 38400 ns,
	      "0001" after 38600 ns,
	      "0010" after 38800 ns,
	      "0011" after 39000 ns,
	      "0100" after 39200 ns,
	      "0101" after 39400 ns,
	      "0110" after 39600 ns,
	      "0111" after 39800 ns,
	      "1000" after 40000 ns,
	      "1001" after 40200 ns,
	      "1010" after 40400 ns,
	      "1011" after 40600 ns,
	      "1100" after 40800 ns,
	      "1101" after 41000 ns,
	      "1110" after 41200 ns,
	      "1111" after 41400 ns,
              --1101
              "0000" after 41600 ns,
	      "0001" after 41800 ns,
	      "0010" after 42000 ns,
	      "0011" after 42200 ns,
	      "0100" after 42400 ns,
	      "0101" after 42600 ns,
	      "0110" after 42800 ns,
	      "0111" after 43000 ns,
	      "1000" after 43200 ns,
	      "1001" after 43400 ns,
	      "1010" after 43600 ns,
	      "1011" after 43800 ns,
	      "1100" after 44000 ns,
	      "1101" after 44200 ns,
	      "1110" after 44400 ns,
	      "1111" after 44600 ns,
              --1110
              "0000" after 44800 ns,
	      "0001" after 45000 ns,
	      "0010" after 45200 ns,
	      "0011" after 45400 ns,
	      "0100" after 45600 ns,
	      "0101" after 45800 ns,
	      "0110" after 46000 ns,
	      "0111" after 46200 ns,
	      "1000" after 46400 ns,
	      "1001" after 46600 ns,
	      "1010" after 46800 ns,
	      "1011" after 47000 ns,
	      "1100" after 47200 ns,
	      "1101" after 47400 ns,
	      "1110" after 47600 ns,
	      "1111" after 47800 ns,
              --1111
              "0000" after 48000 ns,
	      "0001" after 48200 ns,
	      "0010" after 48400 ns,
	      "0011" after 48600 ns,
	      "0100" after 48800 ns,
	      "0101" after 49000 ns,
	      "0110" after 49200 ns,
	      "0111" after 49400 ns,
	      "1000" after 49600 ns,
	      "1001" after 49800 ns,
	      "1010" after 50000 ns,
	      "1011" after 50200 ns,
	      "1100" after 50400 ns,
	      "1101" after 50600 ns,
	      "1110" after 50800 ns,
	      "1111" after 51000 ns;
              


    DUT: entity work.bitComparator
    port map(
      a => a_tb,
      b => b_tb,
      sig => '0',
      lg =>  lg_tb,
      eq => eq_tb,
      ls => ls_tb
    );
end architecture testbench;
